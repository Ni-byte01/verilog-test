`timescale 1ns/1ns
module xor_gate_df(input a,b, output y);
   assign y= a ^ b;
endmodule