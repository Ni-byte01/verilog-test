`timescale 1ns/1ns
module or_gate_df(input a,b, output y);
   assign y= a | b;
endmodule